interface gold_wrapper_if(clk);
input clk;
bit MOSI, SS_n,  rst_n;
bit MISO;
endinterface